/*
Copyright by Nicola Nicolici
Department of Electrical and Computer Engineering
McMaster University
Ontario, Canada
*/

class scoreboard;
   
	mailbox mon2scb;
  
	function new(mailbox mon2scb);
		this.mon2scb = mon2scb;
	endfunction
  
	task main();
	endtask
  
endclass
